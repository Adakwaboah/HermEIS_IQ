library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
-- use IEEE.STD_LOGIC_ARITH.ALL;
-- use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity SineWaveGenerator is
    generic(
        dds_bits :  natural := 32;
        freq_bits:  natural := 32--(dds_bit-log2(100M) + log2(100k));
    );
    Port (
        clk         : in STD_LOGIC;
        reset       : in STD_LOGIC;
        sine_out    : out STD_LOGIC_VECTOR(9 downto 0); -- 10-bit output (adjust size as needed)
        freq_out    : in  std_logic_vector(freq_bits-1 downto 0)
        );
end SineWaveGenerator;

architecture Behavioral of SineWaveGenerator is
    constant TABLE_SIZE : integer := 1024; -- Number of elements in the lookup table
    constant TABLE_WIDTH : integer := 10;   -- Width of each table entry (adjust as needed)
    -- constant fcw_scalar  :  integer := integer(real(2**32/100_000_000));
    constant fcw_scalar  :  integer := integer(real(2**32/(2**26)));
    
    type sine_table_type is array (0 to TABLE_SIZE-1) of STD_LOGIC_VECTOR(TABLE_WIDTH-1 downto 0);


    constant sine_table : sine_table_type :=(
        "1000000000", "1000000011", "1000000110", "1000001001", "1000001100", "1000001111", "1000010010", "1000010101", 
        "1000011001", "1000011100", "1000011111", "1000100010", "1000100101", "1000101000", "1000101011", "1000101111", 
        "1000110010", "1000110101", "1000111000", "1000111011", "1000111110", "1001000001", "1001000100", "1001000111", 
        "1001001011", "1001001110", "1001010001", "1001010100", "1001010111", "1001011010", "1001011101", "1001100000", 
        "1001100011", "1001100110", "1001101001", "1001101101", "1001110000", "1001110011", "1001110110", "1001111001", 
        "1001111100", "1001111111", "1010000010", "1010000101", "1010001000", "1010001011", "1010001110", "1010010001", 
        "1010010100", "1010010111", "1010011010", "1010011101", "1010100000", "1010100011", "1010100110", "1010101001", 
        "1010101100", "1010101111", "1010110010", "1010110101", "1010111000", "1010111011", "1010111101", "1011000000", 
        "1011000011", "1011000110", "1011001001", "1011001100", "1011001111", "1011010010", "1011010101", "1011010111", 
        "1011011010", "1011011101", "1011100000", "1011100011", "1011100101", "1011101000", "1011101011", "1011101110", 
        "1011110001", "1011110011", "1011110110", "1011111001", "1011111100", "1011111110", "1100000001", "1100000100", 
        "1100000110", "1100001001", "1100001100", "1100001110", "1100010001", "1100010100", "1100010110", "1100011001", 
        "1100011100", "1100011110", "1100100001", "1100100011", "1100100110", "1100101001", "1100101011", "1100101110", 
        "1100110000", "1100110011", "1100110101", "1100111000", "1100111010", "1100111101", "1100111111", "1101000010", 
        "1101000100", "1101000110", "1101001001", "1101001011", "1101001110", "1101010000", "1101010010", "1101010101", 
        "1101010111", "1101011001", "1101011100", "1101011110", "1101100000", "1101100010", "1101100101", "1101100111", 
        "1101101001", "1101101011", "1101101110", "1101110000", "1101110010", "1101110100", "1101110110", "1101111000", 
        "1101111010", "1101111101", "1101111111", "1110000001", "1110000011", "1110000101", "1110000111", "1110001001", 
        "1110001011", "1110001101", "1110001111", "1110010001", "1110010011", "1110010101", "1110010111", "1110011000", 
        "1110011010", "1110011100", "1110011110", "1110100000", "1110100010", "1110100011", "1110100101", "1110100111", 
        "1110101001", "1110101011", "1110101100", "1110101110", "1110110000", "1110110001", "1110110011", "1110110101", 
        "1110110110", "1110111000", "1110111001", "1110111011", "1110111101", "1110111110", "1111000000", "1111000001", 
        "1111000011", "1111000100", "1111000110", "1111000111", "1111001000", "1111001010", "1111001011", "1111001101", 
        "1111001110", "1111001111", "1111010001", "1111010010", "1111010011", "1111010100", "1111010110", "1111010111", 
        "1111011000", "1111011001", "1111011010", "1111011100", "1111011101", "1111011110", "1111011111", "1111100000", 
        "1111100001", "1111100010", "1111100011", "1111100100", "1111100101", "1111100110", "1111100111", "1111101000", 
        "1111101001", "1111101010", "1111101011", "1111101100", "1111101100", "1111101101", "1111101110", "1111101111", 
        "1111110000", "1111110000", "1111110001", "1111110010", "1111110011", "1111110011", "1111110100", "1111110101", 
        "1111110101", "1111110110", "1111110110", "1111110111", "1111110111", "1111111000", "1111111001", "1111111001", 
        "1111111001", "1111111010", "1111111010", "1111111011", "1111111011", "1111111100", "1111111100", "1111111100", 
        "1111111101", "1111111101", "1111111101", "1111111101", "1111111110", "1111111110", "1111111110", "1111111110", 
        "1111111110", "1111111111", "1111111111", "1111111111", "1111111111", "1111111111", "1111111111", "1111111111", 
        "1111111111", "1111111111", "1111111111", "1111111111", "1111111111", "1111111111", "1111111111", "1111111111", 
        "1111111110", "1111111110", "1111111110", "1111111110", "1111111110", "1111111101", "1111111101", "1111111101", 
        "1111111101", "1111111100", "1111111100", "1111111100", "1111111011", "1111111011", "1111111010", "1111111010", 
        "1111111001", "1111111001", "1111111001", "1111111000", "1111110111", "1111110111", "1111110110", "1111110110", 
        "1111110101", "1111110101", "1111110100", "1111110011", "1111110011", "1111110010", "1111110001", "1111110000", 
        "1111110000", "1111101111", "1111101110", "1111101101", "1111101100", "1111101100", "1111101011", "1111101010", 
        "1111101001", "1111101000", "1111100111", "1111100110", "1111100101", "1111100100", "1111100011", "1111100010", 
        "1111100001", "1111100000", "1111011111", "1111011110", "1111011101", "1111011100", "1111011010", "1111011001", 
        "1111011000", "1111010111", "1111010110", "1111010100", "1111010011", "1111010010", "1111010001", "1111001111", 
        "1111001110", "1111001101", "1111001011", "1111001010", "1111001000", "1111000111", "1111000110", "1111000100", 
        "1111000011", "1111000001", "1111000000", "1110111110", "1110111101", "1110111011", "1110111001", "1110111000", 
        "1110110110", "1110110101", "1110110011", "1110110001", "1110110000", "1110101110", "1110101100", "1110101011", 
        "1110101001", "1110100111", "1110100101", "1110100011", "1110100010", "1110100000", "1110011110", "1110011100", 
        "1110011010", "1110011000", "1110010111", "1110010101", "1110010011", "1110010001", "1110001111", "1110001101", 
        "1110001011", "1110001001", "1110000111", "1110000101", "1110000011", "1110000001", "1101111111", "1101111101", 
        "1101111010", "1101111000", "1101110110", "1101110100", "1101110010", "1101110000", "1101101110", "1101101011", 
        "1101101001", "1101100111", "1101100101", "1101100010", "1101100000", "1101011110", "1101011100", "1101011001", 
        "1101010111", "1101010101", "1101010010", "1101010000", "1101001110", "1101001011", "1101001001", "1101000110", 
        "1101000100", "1101000010", "1100111111", "1100111101", "1100111010", "1100111000", "1100110101", "1100110011", 
        "1100110000", "1100101110", "1100101011", "1100101001", "1100100110", "1100100011", "1100100001", "1100011110", 
        "1100011100", "1100011001", "1100010110", "1100010100", "1100010001", "1100001110", "1100001100", "1100001001", 
        "1100000110", "1100000100", "1100000001", "1011111110", "1011111100", "1011111001", "1011110110", "1011110011", 
        "1011110001", "1011101110", "1011101011", "1011101000", "1011100101", "1011100011", "1011100000", "1011011101", 
        "1011011010", "1011010111", "1011010101", "1011010010", "1011001111", "1011001100", "1011001001", "1011000110", 
        "1011000011", "1011000000", "1010111101", "1010111011", "1010111000", "1010110101", "1010110010", "1010101111", 
        "1010101100", "1010101001", "1010100110", "1010100011", "1010100000", "1010011101", "1010011010", "1010010111", 
        "1010010100", "1010010001", "1010001110", "1010001011", "1010001000", "1010000101", "1010000010", "1001111111", 
        "1001111100", "1001111001", "1001110110", "1001110011", "1001110000", "1001101101", "1001101001", "1001100110", 
        "1001100011", "1001100000", "1001011101", "1001011010", "1001010111", "1001010100", "1001010001", "1001001110", 
        "1001001011", "1001000111", "1001000100", "1001000001", "1000111110", "1000111011", "1000111000", "1000110101", 
        "1000110010", "1000101111", "1000101011", "1000101000", "1000100101", "1000100010", "1000011111", "1000011100", 
        "1000011001", "1000010101", "1000010010", "1000001111", "1000001100", "1000001001", "1000000110", "1000000011", 
        "1000000000", "0111111100", "0111111001", "0111110110", "0111110011", "0111110000", "0111101101", "0111101010", 
        "0111100110", "0111100011", "0111100000", "0111011101", "0111011010", "0111010111", "0111010100", "0111010000", 
        "0111001101", "0111001010", "0111000111", "0111000100", "0111000001", "0110111110", "0110111011", "0110111000", 
        "0110110100", "0110110001", "0110101110", "0110101011", "0110101000", "0110100101", "0110100010", "0110011111", 
        "0110011100", "0110011001", "0110010110", "0110010010", "0110001111", "0110001100", "0110001001", "0110000110", 
        "0110000011", "0110000000", "0101111101", "0101111010", "0101110111", "0101110100", "0101110001", "0101101110", 
        "0101101011", "0101101000", "0101100101", "0101100010", "0101011111", "0101011100", "0101011001", "0101010110", 
        "0101010011", "0101010000", "0101001101", "0101001010", "0101000111", "0101000100", "0101000010", "0100111111", 
        "0100111100", "0100111001", "0100110110", "0100110011", "0100110000", "0100101101", "0100101010", "0100101000", 
        "0100100101", "0100100010", "0100011111", "0100011100", "0100011010", "0100010111", "0100010100", "0100010001", 
        "0100001110", "0100001100", "0100001001", "0100000110", "0100000011", "0100000001", "0011111110", "0011111011", 
        "0011111001", "0011110110", "0011110011", "0011110001", "0011101110", "0011101011", "0011101001", "0011100110", 
        "0011100011", "0011100001", "0011011110", "0011011100", "0011011001", "0011010110", "0011010100", "0011010001", 
        "0011001111", "0011001100", "0011001010", "0011000111", "0011000101", "0011000010", "0011000000", "0010111101", 
        "0010111011", "0010111001", "0010110110", "0010110100", "0010110001", "0010101111", "0010101101", "0010101010", 
        "0010101000", "0010100110", "0010100011", "0010100001", "0010011111", "0010011101", "0010011010", "0010011000", 
        "0010010110", "0010010100", "0010010001", "0010001111", "0010001101", "0010001011", "0010001001", "0010000111", 
        "0010000101", "0010000010", "0010000000", "0001111110", "0001111100", "0001111010", "0001111000", "0001110110", 
        "0001110100", "0001110010", "0001110000", "0001101110", "0001101100", "0001101010", "0001101000", "0001100111", 
        "0001100101", "0001100011", "0001100001", "0001011111", "0001011101", "0001011100", "0001011010", "0001011000", 
        "0001010110", "0001010100", "0001010011", "0001010001", "0001001111", "0001001110", "0001001100", "0001001010", 
        "0001001001", "0001000111", "0001000110", "0001000100", "0001000010", "0001000001", "0000111111", "0000111110", 
        "0000111100", "0000111011", "0000111001", "0000111000", "0000110111", "0000110101", "0000110100", "0000110010", 
        "0000110001", "0000110000", "0000101110", "0000101101", "0000101100", "0000101011", "0000101001", "0000101000", 
        "0000100111", "0000100110", "0000100101", "0000100011", "0000100010", "0000100001", "0000100000", "0000011111", 
        "0000011110", "0000011101", "0000011100", "0000011011", "0000011010", "0000011001", "0000011000", "0000010111", 
        "0000010110", "0000010101", "0000010100", "0000010011", "0000010011", "0000010010", "0000010001", "0000010000", 
        "0000001111", "0000001111", "0000001110", "0000001101", "0000001100", "0000001100", "0000001011", "0000001010", 
        "0000001010", "0000001001", "0000001001", "0000001000", "0000001000", "0000000111", "0000000110", "0000000110", 
        "0000000110", "0000000101", "0000000101", "0000000100", "0000000100", "0000000011", "0000000011", "0000000011", 
        "0000000010", "0000000010", "0000000010", "0000000010", "0000000001", "0000000001", "0000000001", "0000000001", 
        "0000000001", "0000000000", "0000000000", "0000000000", "0000000000", "0000000000", "0000000000", "0000000000", 
        "0000000000", "0000000000", "0000000000", "0000000000", "0000000000", "0000000000", "0000000000", "0000000000", 
        "0000000001", "0000000001", "0000000001", "0000000001", "0000000001", "0000000010", "0000000010", "0000000010", 
        "0000000010", "0000000011", "0000000011", "0000000011", "0000000100", "0000000100", "0000000101", "0000000101", 
        "0000000110", "0000000110", "0000000110", "0000000111", "0000001000", "0000001000", "0000001001", "0000001001", 
        "0000001010", "0000001010", "0000001011", "0000001100", "0000001100", "0000001101", "0000001110", "0000001111", 
        "0000001111", "0000010000", "0000010001", "0000010010", "0000010011", "0000010011", "0000010100", "0000010101", 
        "0000010110", "0000010111", "0000011000", "0000011001", "0000011010", "0000011011", "0000011100", "0000011101", 
        "0000011110", "0000011111", "0000100000", "0000100001", "0000100010", "0000100011", "0000100101", "0000100110", 
        "0000100111", "0000101000", "0000101001", "0000101011", "0000101100", "0000101101", "0000101110", "0000110000", 
        "0000110001", "0000110010", "0000110100", "0000110101", "0000110111", "0000111000", "0000111001", "0000111011", 
        "0000111100", "0000111110", "0000111111", "0001000001", "0001000010", "0001000100", "0001000110", "0001000111", 
        "0001001001", "0001001010", "0001001100", "0001001110", "0001001111", "0001010001", "0001010011", "0001010100", 
        "0001010110", "0001011000", "0001011010", "0001011100", "0001011101", "0001011111", "0001100001", "0001100011", 
        "0001100101", "0001100111", "0001101000", "0001101010", "0001101100", "0001101110", "0001110000", "0001110010", 
        "0001110100", "0001110110", "0001111000", "0001111010", "0001111100", "0001111110", "0010000000", "0010000010", 
        "0010000101", "0010000111", "0010001001", "0010001011", "0010001101", "0010001111", "0010010001", "0010010100", 
        "0010010110", "0010011000", "0010011010", "0010011101", "0010011111", "0010100001", "0010100011", "0010100110", 
        "0010101000", "0010101010", "0010101101", "0010101111", "0010110001", "0010110100", "0010110110", "0010111001", 
        "0010111011", "0010111101", "0011000000", "0011000010", "0011000101", "0011000111", "0011001010", "0011001100", 
        "0011001111", "0011010001", "0011010100", "0011010110", "0011011001", "0011011100", "0011011110", "0011100001", 
        "0011100011", "0011100110", "0011101001", "0011101011", "0011101110", "0011110001", "0011110011", "0011110110", 
        "0011111001", "0011111011", "0011111110", "0100000001", "0100000011", "0100000110", "0100001001", "0100001100", 
        "0100001110", "0100010001", "0100010100", "0100010111", "0100011010", "0100011100", "0100011111", "0100100010", 
        "0100100101", "0100101000", "0100101010", "0100101101", "0100110000", "0100110011", "0100110110", "0100111001", 
        "0100111100", "0100111111", "0101000010", "0101000100", "0101000111", "0101001010", "0101001101", "0101010000", 
        "0101010011", "0101010110", "0101011001", "0101011100", "0101011111", "0101100010", "0101100101", "0101101000", 
        "0101101011", "0101101110", "0101110001", "0101110100", "0101110111", "0101111010", "0101111101", "0110000000", 
        "0110000011", "0110000110", "0110001001", "0110001100", "0110001111", "0110010010", "0110010110", "0110011001", 
        "0110011100", "0110011111", "0110100010", "0110100101", "0110101000", "0110101011", "0110101110", "0110110001", 
        "0110110100", "0110111000", "0110111011", "0110111110", "0111000001", "0111000100", "0111000111", "0111001010", 
        "0111001101", "0111010000", "0111010100", "0111010111", "0111011010", "0111011101", "0111100000", "0111100011", 
        "0111100110", "0111101010", "0111101101", "0111110000", "0111110011", "0111110110", "0111111001", "0111111100"

    );
    
    -- signal phase_accumulator : integer range 0 to TABLE_SIZE-1 := 0;
    signal phase_accumulator : unsigned(freq_bits-1 downto 0);
    signal phase_inc : unsigned(freq_bits-1 downto 0);

begin
    

    process(clk, reset)
        variable phase_increment    :   unsigned(freq_bits-1 downto 0);
        variable current_phase      :   unsigned(TABLE_WIDTH-1 downto 0);
    begin
        phase_inc <= phase_increment;
        if reset = '1' then
            phase_accumulator <= (others=>'0');
            sine_out <= (others => '0');
        elsif rising_edge(clk) then
            -- Increment phase accumulator based on frequency of the sine wave
            -- For example, for a 1 Hz sine wave, you can use: phase_accumulator <= phase_accumulator + 1;
            -- For higher frequencies, you can use fractional increments to get more resolution.
            phase_increment := to_unsigned( fcw_scalar * to_integer(unsigned(freq_out)) , freq_bits); --* to_integer(unsigned(freq_out));
            phase_accumulator <= phase_accumulator + phase_increment;
            current_phase := phase_accumulator(freq_bits-1 downto freq_bits-TABLE_WIDTH);
            --phase_accumulator <= (phase_accumulator + 1) mod TABLE_SIZE;
            -- Output the corresponding sine value from the lookup table
            sine_out <= sine_table(to_integer(current_phase));
        end if;
    end process;

end Behavioral;
